class StressAppExecutor extends cdnChiUvmSequence;
endclass
